`timescale 1ns / 1ps



module mux8by1_tb();
wire y;
reg [2:0] s;
reg [7:0] a;
muxusingmux uut(a,s,y);
initial
 begin
 a=8'b10101101;s[1]=0;s[0]=0;s[2]=0;#10;
 a=8'b10101101;s[1]=0;s[0]=1;s[2]=0;#10;
 a=8'b10101101;s[1]=1;s[0]=0;s[2]=0;#10;
 a=8'b10101101;s[1]=1;s[0]=1;s[2]=0;#10;
 a=8'b10101101;s[1]=0;s[0]=0;s[2]=1;#10;
 a=8'b10101101;s[1]=0;s[0]=1;s[2]=1;#10;
 a=8'b10101101;s[1]=1;s[0]=0;s[2]=1;#10;
 a=8'b10101101;s[1]=1;s[0]=1;s[2]=1;#10;
 end
endmodule
